# ====================================================================
#
#	intel_npe_npemh.cdl
#
#	Intel npe ethernet driver
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Mark Salter <msalter@redhat.com>
# Original data:
# Contributors:
# Date:           2005-02-08
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_INTEL_NPE_NPEMH {
    display       "Intel NPE message handling layer"
    description   "Message handling layer for Intel Network Processors."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_INTEL_NPE_REQUIRED

    define_proc {
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_INTEL_NPE_NPEMH_CFG";
    }

    compile -library=libextras.a                \
	IxNpeMh.c IxNpeMhConfig.c IxNpeMhReceive.c IxNpeMhSend.c \
	IxNpeMhSolicitedCbMgr.c IxNpeMhUnsolicitedCbMgr.c

    cdl_component CYGPKG_DEVS_ETH_INTEL_NPE_NPEMH_OPTIONS {
        display "Intel npe ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_INTEL_NPE_NPEMH_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -DCPU=33 -DXSCALE=33 -DNDEBUG -DIX_COMPONENT_NAME=7 \
			     -I$(PREFIX)/include/osal                          \
			     -I$(PREFIX)/include/osal/modules/bufferMgt        \
			     -I$(PREFIX)/include/osal/modules/ioMem            \
			     -I$(PREFIX)/include/osal/modules/ioMem            \
			     -I$(PREFIX)/include/osal/ecos/core                \
			     -I$(PREFIX)/include/osal/ecos/modules/bufferMgt   \
			     -I$(PREFIX)/include/osal/ecos/modules/ioMem       \
			     -I$(PREFIX)/include/osal/ecos/platforms/ixp400    \
			"}
            description   "
                This option modifies the set of compiler flags for
                building the Intel npe ethernet driver package.
                These flags are used in addition to the set of
                global flags."
        }
    }
}
# EOF intel_npe_eth_drivers.cdl
