# ====================================================================
#
#      flash_moab.cdl
#
#      FLASH memory - Hardware support for boot FLASH on TAMS MOAB
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Nick Garnett <nickg@calivar.com>
## Copyright (C) 2003 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas, hmt, jskov, tdrury, nickg
# Original data:  gthomas
# Contributors:   gthomas
# Date:           2001-02-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_FLASH_POWERPC_MOAB {
    display       "TAMS MOAB FLASH memory support"
    description   "FLASH memory device(s) support for MOAB board"

    parent        CYGPKG_IO_FLASH
    active_if     CYGPKG_IO_FLASH
    requires      CYGPKG_HAL_POWERPC_MOAB
    requires      { CYGSEM_DEVS_FLASH_POWERPC_MOAB_BOOT || CYGSEM_DEVS_FLASH_POWERPC_MOAB_MAIN }

    cdl_component CYGSEM_DEVS_FLASH_POWERPC_MOAB_BOOT {
        display       "Boot FLASH support"
        default_value 0
        no_define
        description   "
            This option enables the drivers for the bootstrap FLASH
            device.  Note: this device is not suitable for the RedBoot
            Flash Image System (FIS)."

        compile       moab_flash.c
    
        # Arguably this should do in the generic package
        # but then there is a logic loop so you can never enable it.
        cdl_interface CYGINT_DEVS_FLASH_ATMEL_AT49XXXX_REQUIRED {
            display   "Generic Atmel AM49XXXX driver required"
        }

        implements    CYGINT_DEVS_FLASH_ATMEL_AT49XXXX_REQUIRED
    }

    cdl_component CYGSEM_DEVS_FLASH_POWERPC_MOAB_MAIN {
        display       "Main (NAND) FLASH support"
        default_value 1
        no_define
        description   "
            This option enables the drivers for the main FLASH
            device.  Note: this device can be used for the RedBoot
            Flash Image System (FIS)."

        compile       moab_nand_flash.c

        # Arguably this should do in the generic package
        # but then there is a logic loop so you can never enable it.
        cdl_interface CYGINT_DEVS_FLASH_TOSHIBA_TC58XXX_REQUIRED {
            display   "Generic Toshiba TC58XXX driver required"
        }

        implements    CYGINT_DEVS_FLASH_TOSHIBA_TC58XXX_REQUIRED
    }
}
