# ====================================================================
#
#      startup.cdl
#
#      Infrastructure startup configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      bartv
# Original data:  bartv,hmt
# Contributors:
# Date:           1999-06-13
#
#####DESCRIPTIONEND####
#
# ====================================================================

# =================================================================
# The following options allow particular compatibility modes to be
# enabled, when they require specialised support from the startup
# process. These can affect the environment in which the program
# runs.
#
# CYGSEM_START_UITRON_COMPATIBILITY enables compatibility with uItron.
# You must configure uItron with the correct tasks, and then enabling this
# option starts the uItron subsystem. It does this by invoking the function
# cyg_uitron_start().
#
# Both these can also be done by the user overriding cyg_user_start(),
# cyg_package_start(), or cyg_prestart(). Refer to the documentation on
# how and when to do this.

cdl_option CYGSEM_START_UITRON_COMPATIBILITY {
    display       "Start uITRON subsystem"
    default_value 0
    requires      CYGPKG_UITRON
    active_if     CYGPKG_UITRON
    description   "
        Generate a call to initialize the
        uITRON compatibility subsystem
        within the system version of cyg_package_start().
        This enables compatibility with uITRON.
        You must configure uITRON with the correct tasks before
        starting the uItron subsystem.
        If this is disabled, and you want to use uITRON,
        you must call cyg_uitron_start() from your own
        cyg_package_start() or cyg_userstart()."
}
