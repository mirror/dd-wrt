# ====================================================================
#
#      hal_mips_ar2316.cdl
#
#      MIPS AR2316 SOC HAL package configuration data
#
# ====================================================================
######ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Atheros Communications, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting the copyright
## holders.
## -------------------------------------------
######ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      adrian
# Contributors:
# Date:           2003-10-18
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MIPS_AR2316 {
    display  "AR2316 Atheros SOC"
    parent        CYGPKG_HAL_MIPS
    requires      { ((CYGHWR_HAL_MIPS_MIPS32_CORE == "4Kc") || \
                       (CYGHWR_HAL_MIPS_MIPS32_CORE == "4Kp"))  \
                  }
    include_dir   cyg/hal
    define_header hal_mips_ar2316.h
    description   "
           The AR2316 HAL package provides generic support for the
	   Atheros AR2316 and AR2313 WiSoC's. It is also necessary
           to select a specific board package."

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_mips_mips32.h>"
    }

    cdl_option CYGNUM_CACHE_WRITETHRU {
	display		"Use writethru cache"
	flavor		data
	default_value	1
	description	"Set to 1 if you want ot use writethru cache"
    }	

    cdl_option CYGPKG_HAL_MIPS_CACHE_DEFINED {
	display		"Use Write through cache"
	flavor		booldata
	calculated	{CYGNUM_CACHE_WRITETHRU == 1 ? 1 : 0}
	description	"This option sets the cache to writethru cache"
    }

    compile       platform.S plf_misc.c ser16c550c.c
}
