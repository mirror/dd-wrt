# ====================================================================
#
#      hal_m68k_m68000.cdl
#
#      M68K/M68000 variant architectural HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================

cdl_package CYGPKG_HAL_M68K_MCF52xx_MCF5272 {
    display         "mcf5272 68k/Coldfire variant HAL"
    parent          CYGPKG_HAL_M68K_MCF52xx
    requires        CYGPKG_HAL_M68K_MCF52xx
    implements      CYGINT_HAL_M68K_VARIANT
    hardware
    include_dir     cyg/hal
    define_header   hal_m68k_mcf52xx_mcf5272.h

    description   "The  mcf5272  68k/Coldfire  variant  HAL  package  provides
                generic support for this  processor architecture.  It is  also
                necessary to select a specific target platform HAL package."

    define_proc {
        puts $::cdl_header "#include <pkgconf/hal_m68k_mcf52xx.h>"
    }

    compile     proc_startup.c proc_arch.S proc_misc.c memcpy.c

}

