# ====================================================================
#
#      hal_mips_pb44.cdl
#
#      MIPS Atheros PB44 board HAL package configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2003 Atheros Communications, Inc.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting the copyright
## holders.
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      adrian
# Original data:  
# Contributors:   
# Date:           2003-10-18
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_HAL_MIPS_PB44_ROUTER {
    display  "PB44 Router Atheros board"
    parent        CYGPKG_HAL_MIPS
    requires      CYGPKG_HAL_MIPS_AR7100
    define_header hal_mips_pb44.h
    include_dir   cyg/hal
    description   "
           The PB44 Router Atheros HAL package provides support for the PB44
	   test board which is based on the AR7100 SOC with 16M flash.  It 
	   should be used when targetting the actual hardware."

    implements    CYGINT_HAL_DEBUG_GDB_STUBS
    implements    CYGINT_HAL_DEBUG_GDB_STUBS_BREAK
    implements    CYGINT_HAL_VIRTUAL_VECTOR_SUPPORT
    implements    CYGINT_HAL_VIRTUAL_VECTOR_COMM_BAUD_SUPPORT

    compile	  plf_flash.c board_misc.c

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_mips_pb44.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_PLATFORM_H <pkgconf/hal_mips_ar7100.h>"
    }

    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        legal_values  {"RAM" "ROM" "ROMRAM"}
        default_value {"RAM"}
	no_define
	define -file system.h CYG_HAL_STARTUP
        description   "Use the RAM version to load the ROM version as bootrom"
    }


    cdl_interface CYGINT_DEVS_FLASH_AR7100_REQUIRED {
        display   "pb44 has AR7100 spi FLASH part fitted"
        description   "This option enables the driver for AR7100 FLASH"
    }

    implements    CYGINT_DEVS_FLASH_AR7100_REQUIRED

    # The "-o file" is a workaround for CR100958 - without it the
    # output file would end up in the source directory under CygWin.
    # n.b. grep does not behave itself under win32
    make -priority 1 {
        <PREFIX>/include/cyg/hal/plf_defs.inc : <PACKAGE>/src/plf_mk_defs.c
        $(CC) $(CFLAGS) $(INCLUDE_PATH) -Wp,-MD,plf_defs.tmp -o plf_mk_defs.tmp -S $<
        fgrep .equ plf_mk_defs.tmp | sed s/#// > $@
        @echo $@ ": \\" > $(notdir $@).deps
        @tail --lines=2 plf_defs.tmp >> $(notdir $@).deps
        @echo >> $(notdir $@).deps
        @rm plf_defs.tmp plf_mk_defs.tmp
    }

    # Real-time clock/counter specifics
    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants."
        flavor        none
    
        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            calculated    1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            calculated    100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
            calculated    { 110000000 / CYGNUM_HAL_RTC_DENOMINATOR }
            description   "
                The count and compare registers of the AR7100 are used
                to drive the eCos kernel RTC. The count register
                increments at the CPU clock speed."
        }
    }

    cdl_component CYGNUM_HAL_BOARD_TYPE {
        display       "board type"
        flavor        data
        default_value {"\"pb44-router\""}
        description   "board type string displayed part of version command"
	}

	cdl_option CYGNUM_CONFIG_PRODUCT_ID {
	display	        "PB44 Product ID value"
	flavor          data
	default_value   131
	description     "PB44 Product ID is 131"
    }

    cdl_option CYGNUM_PLL_FREQ {
        display       "PLL config for CPU/DDR/AHB frequencies"
        flavor        data
        calculated    {"AR7100_PLL_680_340_170"}
        description   "PLL config for CPU/DDR/AHB frequencies"
    }

# Number is value to use in ar7100_pll <n> command
#
# AR7100_PLL_USE_REV_ID    0
# AR7100_PLL_200_200_100   1
# AR7100_PLL_300_300_150   2
# AR7100_PLL_333_333_166   3
# AR7100_PLL_266_266_133   4
# AR7100_PLL_266_266_66    5
# AR7100_PLL_400_400_200   6
# AR7100_PLL_600_300_150   7
# AR7100_PLL_680_340_170   8
# AR7100_PLL_720_360_180   30
# AR7100_PLL_800_400_200   31


    cdl_option CYGNUM_CONFIG_SEC_PLL {
	display	        "PLL Secondary Configuration"
	flavor          data
	default_value   0x000050C0
	description     "Initial values for secondary configuration options such as Eth and PCI clocks"
    }
#	default_value   0x000050C0 <--- internal PCI clock */
#	default_value   0x004050C0 <--- external PCI clock */

    cdl_option CYGNUM_CONFIG_ETH_EXT_CLOCK {
	display	        "PLL Configuration Ethernet clock"
	flavor          data
	default_value   0x00001313
	description     "Initial values for PLL Ethernet clock (25MHz)"
    }

    cdl_option CYGNUM_CONFIG_PCI_CLOCK {
	display	        "PLL Configuration PCI clock"
	flavor          data
	default_value   0x000000ee
	description     "Initial values for internal PCI Clock"
    }
#	default_value   0x000000ee <---- 33 MHz
#	default_value   0x00000067 <---- 66 MHz

    cdl_option CYGNUM_RAM_ENTRY {
	display		"Linked entry address"
	flavor		data
	default_value	0x80010000
	description	"Text segment load address."
    }
 
    cdl_option CYGNUM_RAM_SIZE {
        display         "RAM Memory size"
        flavor          data
        default_value   0x2000000
        description     "RAM memory size"
    }

    cdl_option CYGNUM_DDR_REFRESH_VAL {
        display         "DDR Refresh value"
        flavor          data
        default_value   0x461b
        description     "DDR Refresh value"
    }

    cdl_option CYGNUM_DDR_MODE_VAL {
          display         "DDR Mode value"
          flavor          data
          default_value   0x63  
          description     "DDR Mode value, note: startup will change CAS 2.5 -> 3 if DDR >= 400 to 0x33"
    }

    cdl_option CYGNUM_DDR_RD_DATA_THIS_CYCLE_VAL {
          display         "DDR_RD_DATA_THIS_CYCLE value"
          flavor          data
          default_value   0xff
          description     "DDR Read Data This Cycle value "
    }

    cdl_option CYGNUM_DDR_CONFIG_VAL {
          display         "DDR CONFIG value"
          flavor          data
          default_value   0x6fb8884e  
          description     "DDR CONFIG value, note: startup will change CAS 2.5 -> 3 if DDR 400 (0x77b8884e)"
    }

    cdl_option CYGNUM_DDR_CONFIG2_VAL {
          display         "DDR CONFIG2 value"
          flavor          data
          default_value   0x812cd6a8
          description     "DDR CONFIG2 value"
    }

    cdl_option CYGNUM_EFFECTIVE_RAM_SIZE {
        display         "Effective RAM Memory size"
        flavor          data
        calculated      {CYGNUM_RAM_SIZE - 0x10000}
        description     "Effective RAM memory size"
    }

    cdl_option CYGNUM_FLASH_BLOCK_NUM {
        display         "Number of flash blocks"
        flavor          data
        default_value   0x100
        description     "Number of blocks in flash memory"
    }

    cdl_option CYGNUM_FLASH_BLOCK_SIZE {
	display		"Flash block size"
	flavor		data
	default_value	0x10000
	description	"Block size for erasing flash"
    }

    cdl_option CYGNUM_FLASH_SIZE {
	display		"Flash Memory size"
	flavor		data
	calculated	{CYGNUM_FLASH_BLOCK_SIZE * CYGNUM_FLASH_BLOCK_NUM}
	description	"Flash memory size used for memory layout"
    }

    cdl_option CYGNUM_FLASH_BASE {
	display		"Flash base address"
	flavor		data
	default_value	0xbf000000
	description	"Flash BaseAddress for access"
    }

    cdl_option CYGNUM_FLASH_WIDTH {
	display		"Bus width of flash"
	flavor		data
	default_value	16
	description	"Flash memory bus width"
    }

    cdl_option CYGNUM_FLASH_16AS8 {
	flavor		booldata
	default_value	{ CYGNUM_FLASH_WIDTH == 8 ? 1 : 0 }
    }

    cdl_option CYGNUM_FLASH_END_RESERVED_BYTES {
	display		"Reserved room at end of flash"
	flavor		data
	calculated	0x10000
	description	"Important information is placed at the end of flash
		         by the manufacturer.  It must not be modified or
			 erased, or the board may not function correctly."
    }

    cdl_option CYGNUM_INIT_SP_OFFSET {
	display		"Temporary init stack offset"
	flavor		data
	default_value	0x1000
	description	"Base for temp stack used during init"
    }

    cdl_option CYGNUM_USE_ENET_PHY {
        display		"Selects which enet phy to use"
        flavor          data
        default_value   {AR7100_VSC8601_ENET_PHY}
        description	"PHY configuration for MAC0/1"
    }

    cdl_option CYGNUM_GE0_IFTYPE {
        display		"Selects interface type on GE port 0"
        flavor          data
        calculated      {"AR7100_IF_RGMII"}
        description	"RGMII interface on port 0"
    }

    cdl_option CYGNUM_GE1_IFTYPE {
        display		"Selects interface type on GE port 1"
        flavor          data
        calculated      {"AR7100_IF_RGMII"}
        description	"RGMII interface on port 1"
    }

    cdl_option CYGBLD_BUILD_GDB_STUBS {
	display "Build GDB stub ROM image"
	default_value 0
	parent CYGBLD_GLOBAL_OPTIONS
	requires { CYG_HAL_STARTUP == "ROM" }
	requires CYGSEM_HAL_ROM_MONITOR
	requires CYGBLD_BUILD_COMMON_GDB_STUBS
	requires CYGDBG_HAL_DEBUG_GDB_INCLUDE_STUBS
	requires ! CYGDBG_HAL_DEBUG_GDB_BREAK_SUPPORT
	requires ! CYGDBG_HAL_DEBUG_GDB_THREAD_SUPPORT
	requires ! CYGDBG_HAL_COMMON_INTERRUPTS_SAVE_MINIMUM_CONTEXT
	requires ! CYGDBG_HAL_COMMON_CONTEXT_SAVE_MINIMUM
	no_define
	description "
                This option enables the building of the GDB stubs for the
                board. The common HAL controls takes care of most of the
                build process, but the final conversion from ELF image to
                binary data is handled by the platform CDL, allowing
                relocation of the data if necessary."

	make -priority 320 {
	    <PREFIX>/bin/gdb_module.bin : <PREFIX>/bin/gdb_module.img
	    $(OBJCOPY) -O binary $< $@
	}
    }

    cdl_option CYGNUM_HAL_BREAKPOINT_LIST_SIZE {
        display       "Number of breakpoints supported by the HAL."
        flavor        data
        default_value 25
        description   "
            This option determines the number of breakpoints supported by the HAL."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display      "Number of communication channels on the board"
        flavor       data
        calculated   1
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The AR7100 has only one serial port. This option
           chooses which port will be used to connect to a host
           running GDB."
    }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
        display          "Diagnostic serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    0
        description      "
           The AR7100 has only one serial port.  This option
           chooses which port will be used for diagnostic output."
     }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CHANNELS_DEFAULT_BAUD {
        display       "Console/GDB serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        define        CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD
        description   "
            This option controls the default baud rate used for the
            Console/GDB connection."
    }

    cdl_component CYGHWR_MEMORY_LAYOUT {
        display "Memory layout"
        flavor data
        no_define
        calculated { CYG_HAL_STARTUP == "RAM" ? "mips_pb44_ram" : \
                     CYG_HAL_STARTUP == "ROMRAM" ? "mips_pb44_romram" : \
                                                "mips_pb44_rom" }

        cdl_option CYGHWR_MEMORY_LAYOUT_LDI {
            display "Memory layout linker script fragment"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_LDI
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_mips_pb44_ram.ldi>" : \
                         CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_mips_pb44_romram.ldi>" : \
                                                    "<pkgconf/mlt_mips_pb44_rom.ldi>" }
        }

        cdl_option CYGHWR_MEMORY_LAYOUT_H {
            display "Memory layout header file"
            flavor data
            no_define
            define -file system.h CYGHWR_MEMORY_LAYOUT_H
            calculated { CYG_HAL_STARTUP == "RAM" ? "<pkgconf/mlt_mips_pb44_ram.h>" : \
                         CYG_HAL_STARTUP == "ROMRAM" ? "<pkgconf/mlt_mips_pb44_romram.h>" : \
                                                    "<pkgconf/mlt_mips_pb44_rom.h>" }
        }
    }

    cdl_option CYGSEM_HAL_USE_ROM_MONITOR {
        display       "Work with a ROM monitor"
        flavor        booldata
        legal_values  { "Generic" "GDB_stubs" }
        default_value { CYG_HAL_STARTUP == "RAM" ? "GDB_stubs" : 0 }
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { CYG_HAL_STARTUP == "RAM" }
        description   "
            Support can be enabled for three different varieties of ROM monitor.
            This support changes various eCos semantics such as the encoding
            of diagnostic output, or the overriding of hardware interrupt
            vectors.
            Firstly there is \"Generic\" support which prevents the HAL
            from overriding the hardware vectors that it does not use, to
            instead allow an installed ROM monitor to handle them. This is
            the most basic support which is likely to be common to most
            implementations of ROM monitor.
            \"GDB_stubs\" provides support when GDB stubs are
            included in the ROM monitor or boot ROM."
    }

    cdl_option CYGSEM_HAL_ROM_MONITOR {
        display       "Behave as a ROM monitor"
        flavor        bool
        default_value 0
        parent        CYGPKG_HAL_ROM_MONITOR
        requires      { (CYG_HAL_STARTUP == "ROM") || (CYG_HAL_STARTUP == "ROMRAM") }
        description   "
            Enable this option if this program is to be used as a ROM monitor,
            i.e. applications will be loaded into RAM on the board, and this
            ROM monitor may process exceptions or interrupts generated from the
            application. This enables features such as utilizing a separate
            interrupt stack when exceptions are generated."
    }

    cdl_component CYGPKG_CYGMON_HAL_OPTIONS {
        display       "CygMon HAL options"
        flavor        none
        no_define
        parent        CYGPKG_CYGMON
        active_if     CYGPKG_CYGMON
        description   "
            This option also lists the target's requirements for a valid CygMon
            configuration."

        cdl_option CYGBLD_BUILD_CYGMON_BIN {
            display       "Build CygMon ROM binary image"
            active_if     CYGBLD_BUILD_CYGMON
            default_value 1
            no_define
            description "This option enables the conversion of the CygMon ELF
                         image to a binary image suitable for ROM programming."
    
            make -priority 325 {
                <PREFIX>/bin/cygmon.srec : <PREFIX>/bin/cygmon.elf
                $(OBJCOPY) --strip-debug $< $(@:.bin=.img) 
                $(OBJCOPY) -O srec $< $@
            }
        }
    }

    cdl_component CYGPKG_REDBOOT_HAL_OPTIONS {
        display       "Redboot HAL options"
        flavor        none
        no_define
        parent        CYGPKG_REDBOOT
        active_if     CYGPKG_REDBOOT
        description   "
            This option lists the target's requirements for a valid Redboot
            configuration."

        cdl_option CYGBLD_BUILD_REDBOOT_BIN {
            display       "Build Redboot ROM binary image"
            active_if     CYGBLD_BUILD_REDBOOT
            default_value 1
            no_define
            description "This option enables the conversion of the Redboot ELF
                         image to a binary image suitable for ROM programming."
    
            compile -library=libextras.a
    
            make -priority 325 {
                <PREFIX>/bin/redboot.srec : <PREFIX>/bin/redboot.elf
                $(OBJCOPY) --strip-all $< $(@:.srec=.img)
                $(OBJCOPY) -O srec $< $@
            }
        }
    }
}
