# ====================================================================
#
#      cpuload.cdl
#
#      cpu load measurements
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 2002 Andrew Lunn
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Andrew Lunn
# Original data:  Andrew Lunn
# Contributors:
# Date:           2002-08-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_CPULOAD {
    display       "Measure the current CPU load"
    requires      CYGPKG_KERNEL
    requires      !CYGPKG_KERNEL_SMP_SUPPORT
    include_dir   cyg/cpuload
    
    compile cpuload.cxx
    description "
       This package measures the CPU load over the last 100ms, 1second 
       and 10 second. All loads are returned as a percentage, ie 0-100.
       This is only a rough measure. Any clever power management, sleep 
       modes etc, will cause these results to be wrong."
    doc           ref/services-cpuload.html

    cdl_option CYGPKG_CPULOAD_TESTS {
        display "CPU load measurement tests"
        flavor  data   
        no_define      
        calculated { "tests/cpuload" }
    }
}

