#====================================================================
#
#      rattler_eth_drivers.cdl
#
#      Hardware specifics for A&M Rattler ethernet
#
#====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      gthomas, hmt
# Original data:  gthomas
# Contributors:   gthomas, F.Robbins
# Date:           2003-08-19
#
#####DESCRIPTIONEND####
#
#====================================================================

cdl_package CYGPKG_DEVS_ETH_POWERPC_RATTLER {
    display       "A&M Rattler (MPC8250) ethernet support"
    description   "Hardware specifics for A&M Rattler ethernet"

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_IO_ETH_DRIVERS
    active_if	  CYGPKG_HAL_POWERPC 
    active_if	  CYGPKG_HAL_POWERPC_MPC8XXX

    requires      CYGPKG_DEVS_ETH_POWERPC_FCC
    requires      CYGPKG_HAL_POWERPC_RATTLER
    requires      CYGHWR_DEVS_ETH_PHY_AM79C874

    cdl_option CYGHWR_DEVS_ETH_POWERPC_RATTLER_FCC1 {
        display       "Include fcc1/eth0 ethernet device"
        default_value 1
        description   "
          This option controls whether a driver for FCC1/eth0
          is included in the resulting system."
        implements    CYGHWR_NET_DRIVERS
        implements    CYGHWR_NET_DRIVER_ETH0
    }

    cdl_option CYGHWR_DEVS_ETH_POWERPC_RATTLER_FCC2 {
        display       "Include fcc2/eth1 ethernet device"
        default_value 1
        description   "
          This option controls whether a driver for FCC2/eth1
          is included in the resulting system."
        implements    CYGHWR_NET_DRIVERS
        implements    CYGHWR_NET_DRIVER_ETH1
        requires      CYGHWR_DEVS_ETH_POWERPC_RATTLER_FCC1
    }

    include_dir   cyg/io

    define_proc {
        puts $::cdl_system_header "#define CYGDAT_DEVS_FCC_ETH_CDL <pkgconf/devs_eth_powerpc_rattler.h>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_FCC_ETH_INL <cyg/io/rattler_eth.inl>"
    }
}
