# ====================================================================
#
#       ixdp425_npe_eth_driver.cdl
#
#       Ethernet driver
#       IXDP425 and builting NPE support
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter
# Original data:  hmt
# Contributors:   gthomas
# Date:           2003-03-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_ARM_IXDP425_NPE {
    display       "IXDP425 with builtin NPE ethernet driver"
    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_HAL_ARM_XSCALE_IXDP425
    requires      CYGPKG_DEVS_ETH_INTEL_NPE

    include_dir   cyg/io

    # FIXME: This really belongs in the INTEL_NPE package
    cdl_interface CYGINT_DEVS_ETH_INTEL_NPE_REQUIRED {
        display   "Intel Network Processor ethernet driver required"
    }

    define_proc {
        puts $::cdl_system_header "/***** ethernet driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_INTEL_NPE_INL <cyg/io/ixdp425_npe.inl>"
 
 	puts $::cdl_system_header "#define CYGDAT_DEVS_ETH_INTEL_NPE_CFG <pkgconf/devs_eth_arm_ixdp425_npe.h>"

        puts $::cdl_system_header "/*****  ethernet driver proc output end  *****/"
    }


    cdl_component CYGPKG_DEVS_ETH_ARM_IXDP425_NPE_ETH0 {
        display       "IXDP425 ethernet port driver for NPE B"
        flavor        bool
        default_value 1
        description   "
            This option includes the IXDP425 ethernet device driver for
            builtin NPE B."

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH0
        implements CYGINT_DEVS_ETH_INTEL_NPE_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_ARM_IXDP425_NPE_ETH0_NAME {
            display       "Device name for the ETH0 ethernet port driver"
            flavor        data
            default_value {"\"eth0\""}
            description   "
                This option sets the name of the ethernet device for a
                NPEB-based ethernet port."
        }
    }

    cdl_component CYGPKG_DEVS_ETH_ARM_IXDP425_NPE_ETH1 {
        display       "IXDP425 ethernet port driver for NPE C"
        flavor        bool
        default_value 1
        description   "
            This option includes the IXDP425 ethernet device driver for
            builtin NPE C."

        implements CYGHWR_NET_DRIVERS
        implements CYGHWR_NET_DRIVER_ETH1
        implements CYGINT_DEVS_ETH_INTEL_NPE_REQUIRED

        cdl_option CYGDAT_DEVS_ETH_ARM_IXDP425_NPE_ETH1_NAME {
            display       "Device name for the ETH1 ethernet port driver"
            flavor        data
            default_value {"\"eth1\""}
            description   "
                This option sets the name of the ethernet device for a
                NPEC-based ethernet port."
        }
    }

    cdl_option CYGSEM_DEVS_ETH_INTEL_NPE_PLATFORM_EEPROM {
        display       "Platform uses EEPROM to hold MAC addresses."
        flavor bool
        default_value 1
    }
}

