# ====================================================================
#
#	intel_npe_eth_drivers.cdl
#
#	Intel npe ethernet driver
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      msalter, from i82544 original
# Original data:  hmt, nickg
# Contributors:	  hmt, gthomas, jskov
# Date:           2003-03-20
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVS_ETH_INTEL_NPE {
    display       "Intel NPE ethernet driver"
    description   "Ethernet driver for Intel Network Processors."

    parent        CYGPKG_IO_ETH_DRIVERS
    active_if     CYGPKG_IO_ETH_DRIVERS

    active_if     CYGINT_DEVS_ETH_INTEL_NPE_REQUIRED

    define_proc {
        puts $::cdl_header "#include CYGDAT_DEVS_ETH_INTEL_NPE_CFG";
    }

    compile       -library=libextras.a if_npe.c \
	IxOsalOsServices.c IxOsalOsCacheMMU.c IxOsalOsThread.c  \
	IxOsalIoMem.c IxOsalBufferMgt.c \
	IxOsalOsMsgQ.c IxOsalOsSemaphore.c

    cdl_option CYGDBG_DEVS_ETH_INTEL_NPE_CHATTER {
	display "Prints ethernet device status info during startup"
	default_value 0
	description   "
	    The ethernet device initialization code can print lots of info
	    to confirm that it has found the devices, read the MAC address
            from EEPROM correctly, and so on, and also displays the mode
            (10/100MHz, half/full duplex) of the connection."
    }

    cdl_option CYGNUM_DEVS_ETH_INTEL_NPE_DEV_COUNT {
	display "Number of supported interfaces."
	calculated    { CYGINT_DEVS_ETH_INTEL_NPE_REQUIRED }
        flavor        data
	description   "
	    This option selects the number of PCI ethernet interfaces to
            be supported by the driver."
    }

    cdl_option CYGNUM_DEVS_ETH_INTEL_NPE_MAX_RX_DESCRIPTORS {
        display       "Maximum number of RX descriptors"
        flavor  data
        default_value { CYGPKG_REDBOOT ? 4 : 64 }
        define        MAX_RX_DESCRIPTORS
        description   "
                An RX descriptor is used for each ethernet frame required
                to be passed to the upper networking layers. This option
                sets the maximum number of these. Higher numbers use more
                memory, lower numbers will reduce performance. The system
                appears to work OK with as few as 8 descriptors but limps
                painfully with only 4. Performance is better with more than
                8, but assuming the size of non-cached (so useless for anything
                else) memory window is 1Mb, we might as well use it all.
                128 RX and TX descriptors uses the whole 1Mb, near enough."
    }
    
    cdl_option CYGNUM_DEVS_ETH_INTEL_NPE_MAX_TX_DESCRIPTORS {
        display       "Maximum number of TX descriptors"
        flavor  data
        default_value { CYGPKG_REDBOOT ? 2 : 64 }
        define        MAX_TX_DESCRIPTORS
        description   "
                A TX descriptor is used for each ethernet frame passed down
                from upper networking layers for transmission. This option
                sets the maximum number of these. Higher numbers use more
                memory, lower numbers will reduce performance. The system
                appears to work OK with as few as 8 descriptors but limps
                painfully with only 4. Performance is better with more than
                8, but assuming the size of non-cached (so useless for anything
                else) memory window is 1Mb, we might as well use it all.
                128 RX and TX descriptors uses the whole 1Mb, near enough."
    }

    cdl_interface CYGINT_DEVS_ETH_INTEL_NPEA_SMII {
	display "Support SMII PHY on NPE-A"
    }

    cdl_interface CYGINT_DEVS_ETH_INTEL_NPEB_SMII {
	display "Support SMII PHY on NPE-B"
    }

    cdl_interface CYGINT_DEVS_ETH_INTEL_NPEC_SMII {
	display "Support SMII PHY on NPE-C"
    }

    cdl_interface CYGINT_DEVS_ETH_INTEL_NPE_PHY_DISCOVERY {
	display "Support determination of NPE/PHY connection at runtime."
    }

    cdl_component CYGPKG_DEVS_ETH_INTEL_NPE_REDBOOT_HOLDS_UTOPIA_FLAG {
	display         "RedBoot manages flag indicating if UTOPIA on NPE-A"
	flavor          bool
	default_value	1

	active_if     CYGSEM_HAL_VIRTUAL_VECTOR_SUPPORT
	active_if     { CYGHWR_HAL_ARM_XSCALE_CPU == "IXP46x" }

	description   "Enabling this option will allow the UTOPIA flag to be
                       acquired from RedBoot's configuration data, stored in
                       flash memory."

	cdl_component CYGPKG_DEVS_ETH_INTEL_NPE_REDBOOT_HOLDS_UTOPIA_FLAG_VAR {
	    display        "Build-in flash config field for UTOPIA flag"
	    flavor         bool
	    default_value  1

	    active_if       CYGPKG_REDBOOT
	    active_if       CYGPKG_REDBOOT_FLASH
	    active_if       CYGSEM_REDBOOT_FLASH_CONFIG
	    active_if 	    CYGPKG_REDBOOT_NETWORKING

	    description	"
	    This option controls the presence of RedBoot flash
	    configuration fields for the UTOPIA flag when you
	    are building RedBoot. This option cannot be enabled
            outside of building RedBoot."
	}
    }

    cdl_option CYGDAT_DEVS_ETH_INTEL_NPE_DEFAULT_UTOPIA_FLAG {
        display       "The UTOPIA flag default"
        flavor        bool
        default_value 1
	active_if     { CYGHWR_HAL_ARM_XSCALE_CPU == "IXP46x" }
	description	"
	    This option is the default value of the UTOPIA flag. If
            true, NPE-A is used for UTOPIA. If the flag is false,
            NPE-A is used for ethernet. If RedBoot is used to hold
            the UTOPIA flag, this option is used to set the default
            value which may be overridden with the RedBoot fconfig
            command."
    }

    cdl_component CYGPKG_DEVS_ETH_INTEL_NPE_REDBOOT_HOLDS_ESA {
	display         "RedBoot manages ESA data"
	flavor          bool
	default_value	1

	active_if     CYGSEM_HAL_VIRTUAL_VECTOR_SUPPORT
	active_if     !CYGSEM_DEVS_ETH_INTEL_NPE_PLATFORM_EEPROM

	description   "Enabling this option will allow the ethernet
	station address to be acquired from RedBoot's configuration data,
	stored in flash memory.  It can be overridden individually by the
	'Set the ethernet station address' option for each interface."

	cdl_component CYGPKG_DEVS_ETH_INTEL_NPE_REDBOOT_HOLDS_ESA_VARS {
	    display        "Build-in flash config fields for ESAs"
	    flavor         bool
	    default_value  1

	    active_if       CYGPKG_REDBOOT
	    active_if       CYGPKG_REDBOOT_FLASH
	    active_if       CYGSEM_REDBOOT_FLASH_CONFIG
	    active_if 	    CYGPKG_REDBOOT_NETWORKING

	    description	"
	    This option controls the presence of RedBoot flash
	    configuration fields for the ESAs of the interfaces when you
	    are building RedBoot.  It is independent of whether RedBoot
	    itself uses the network or any particular interface."
	}
    }

    cdl_component CYGPKG_DEVS_ETH_INTEL_NPE_OPTIONS {
        display "Intel npe ethernet driver build options"
        flavor  none
	no_define

        cdl_option CYGPKG_DEVS_ETH_INTEL_NPE_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "-D_KERNEL -D__ECOS -DCPU=33 -DXSCALE=33 -DSKIP_NPE_LINK_CHECK           \
                             -DIX_COMPONENT_NAME=1 -DNDEBUG                    \
			     -I$(PREFIX)/include/osal                          \
			     -I$(PREFIX)/include/osal/modules/bufferMgt        \
			     -I$(PREFIX)/include/osal/modules/ioMem            \
			     -I$(PREFIX)/include/osal/modules/ioMem            \
			     -I$(PREFIX)/include/osal/ecos/core                \
			     -I$(PREFIX)/include/osal/ecos/modules/bufferMgt   \
			     -I$(PREFIX)/include/osal/ecos/modules/ioMem       \
			     -I$(PREFIX)/include/osal/ecos/platforms/ixp400    \
			"}
            description   "
                This option modifies the set of compiler flags for
                building the Intel npe ethernet driver package.
                These flags are used in addition to the set of
                global flags."
        }
    }
}
# EOF intel_npe_eth_drivers.cdl
