# ====================================================================
#
#      wallclock_ref4955.cdl
#
#      eCos wallclock for REF4955 driver configuration data
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      jskov
# Contributors:   jskov
# Date:           2000-05-25
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK_MIPS_REF4955 {
    parent        CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_IO_WALLCLOCK
    display       "REF4955 wallclock driver"
    requires      CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1742
    requires      CYGPKG_HAL_MIPS_TX49_REF4955
    hardware
    compile       wallclock_ref4955.cxx
    implements    CYGINT_WALLCLOCK_HW_IMPLEMENTATIONS
    implements    CYGINT_WALLCLOCK_SET_GET_MODE_SUPPORTED
    active_if     CYGIMP_WALLCLOCK_HARDWARE

    cdl_option CYGIMP_WALLCLOCK_HARDWARE {
        parent    CYGPKG_IO_WALLCLOCK_IMPLEMENTATION
        display       "Hardware wallclock"
        default_value 1
        implements    CYGINT_WALLCLOCK_IMPLEMENTATIONS
    }

    cdl_component CYGPKG_DEVICES_WALLCLOCK_MIPS_REF4955_OPTIONS {
        display "REF4955 wallclock build options"
        flavor  none
        description   "
	    Package specific build options including control over
	    compiler flags used only in building this package,
	    and details of which tests are built."


        cdl_option CYGPKG_DEVICES_WALLCLOCK_MIPS_REF4955_CFLAGS_ADD {
            display "Additional compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are used in addition
                to the set of global flags."
        }

        cdl_option CYGPKG_DEVICES_WALLCLOCK_MIPS_REF4955_CFLAGS_REMOVE {
            display "Suppressed compiler flags"
            flavor  data
            no_define
            default_value { "" }
            description   "
                This option modifies the set of compiler flags for
                building the wallclock device. These flags are removed from
                the set of global flags if present."
        }

    }
}
