# ====================================================================
#
#      moab_wallclock_drivers.cdl
#
#      Wallclock drivers - support for DS1307 RTC on the TAMS MOAB
#
# ====================================================================
#####ECOSGPLCOPYRIGHTBEGIN####
## -------------------------------------------
## This file is part of eCos, the Embedded Configurable Operating System.
## Copyright (C) 1998, 1999, 2000, 2001, 2002 Red Hat, Inc.
## Copyright (C) 2003 Gary Thomas
##
## eCos is free software; you can redistribute it and/or modify it under
## the terms of the GNU General Public License as published by the Free
## Software Foundation; either version 2 or (at your option) any later version.
##
## eCos is distributed in the hope that it will be useful, but WITHOUT ANY
## WARRANTY; without even the implied warranty of MERCHANTABILITY or
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License
## for more details.
##
## You should have received a copy of the GNU General Public License along
## with eCos; if not, write to the Free Software Foundation, Inc.,
## 59 Temple Place, Suite 330, Boston, MA 02111-1307 USA.
##
## As a special exception, if other files instantiate templates or use macros
## or inline functions from this file, or you compile this file and link it
## with other works to produce a work based on this file, this file does not
## by itself cause the resulting work to be covered by the GNU General Public
## License. However the source code for this file must still be made available
## in accordance with section (3) of the GNU General Public License.
##
## This exception does not invalidate any other reasons why a work based on
## this file might be covered by the GNU General Public License.
##
## Alternative licenses for eCos may be arranged by contacting Red Hat, Inc.
## at http://sources.redhat.com/ecos/ecos-license/
## -------------------------------------------
#####ECOSGPLCOPYRIGHTEND####
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      rajt
# Contributors:   rajt
# Date:           2001-07-19
#
#####DESCRIPTIONEND####
#
# ====================================================================

cdl_package CYGPKG_DEVICES_WALLCLOCK_POWERPC_MOAB {
    display       "TAMS MOAB board RTC Driver"
    description   "RTC driver for TAMS MOAB."

    parent        CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_IO_WALLCLOCK
    active_if     CYGPKG_HAL_POWERPC_MOAB
    requires      CYGPKG_DEVICES_WALLCLOCK_DALLAS_DS1307

    include_dir   cyg/io

    define_proc {
        puts $::cdl_system_header "/***** MOAB RTC driver proc output start *****/"
        puts $::cdl_system_header "#define CYGDAT_DEVS_WALLCLOCK_DALLAS_1307_INL <cyg/io/devices_wallclock_moab.inl>"
        puts $::cdl_system_header "#define CYGDAT_DEVS_WALLCLOCK_MOAB_CFG <pkgconf/devices_wallclock_powerpc_moab.h>"
        puts $::cdl_system_header "/***** MOAB RTC driver proc output end  *****/"
    }
}
